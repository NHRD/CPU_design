library IEEE;
use IEEE.std_logic_1164.all;

entity adder_4bit is
    port(
        BIN :   in std_logic_vector(3 downto 0);
        SUM :   out std_logic_vector(6 downto 0)
    );
end adder_4bit;

architecture RTL of dec_7seg_hdl is

    signal not_BIN(0)   :   std_logic_vector

begin
    

end RTL;

